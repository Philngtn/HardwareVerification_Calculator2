`include "driver.sv"
`include "generator.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "monitor.sv"
`include "checker.sv"


