library verilog;
use verilog.vl_types.all;
entity checker_sv_unit is
end checker_sv_unit;
