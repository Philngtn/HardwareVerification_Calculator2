library verilog;
use verilog.vl_types.all;
entity environment_sv_unit is
end environment_sv_unit;
