library verilog;
use verilog.vl_types.all;
entity cal_trans_sv_unit is
end cal_trans_sv_unit;
