library verilog;
use verilog.vl_types.all;
entity testDrive_sv_unit is
end testDrive_sv_unit;
