library verilog;
use verilog.vl_types.all;
entity cal_if is
    port(
        clk             : in     vl_logic
    );
end cal_if;
