library verilog;
use verilog.vl_types.all;
entity transaction_sv_unit is
end transaction_sv_unit;
