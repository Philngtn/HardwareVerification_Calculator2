library verilog;
use verilog.vl_types.all;
entity generator_sv_unit is
end generator_sv_unit;
