library verilog;
use verilog.vl_types.all;
entity agent_sv_unit is
end agent_sv_unit;
