library verilog;
use verilog.vl_types.all;
entity cal_ifc_sv_unit is
end cal_ifc_sv_unit;
